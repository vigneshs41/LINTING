module OR2(
  input A, B,
  output Y
);
  assign Y = A | B;
endmodule

